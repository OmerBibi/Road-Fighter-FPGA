//-- feb 2021 add all colors square 
// (c) Technion IIT, Department of Electrical Engineering 2021


module	ROADRGB	(	

					input	logic	clk,
					input	logic	resetN,
					input	logic	startOfFrame,
					input logic	[10:0]	pixelX,
					input logic	[10:0]	pixelY,
					input	logic	InsideRectangle,
					input	logic	[1:0] speed,
					output	logic	[7:0]	BG_RGB,
					output	logic		boardersDrawReq 
);



localparam logic [7:0] BLACK_COLOR = 8'b00000000;
localparam logic [7:0] LIGHT_GRAY_COLOR = 8'b10110110;
localparam logic [7:0] DARK_GRAY_COLOR = 8'b01101101;
localparam logic [7:0] WHITE_COLOR = 8'b11111111;
localparam logic [7:0] SEA_COLOR = 8'b10011011;
localparam logic [7:0] SEA2_COLOR = 8'b01111011;
localparam logic [7:0] SAND_COLOR = 8'b11111101;
localparam logic [7:0] GREEN_COLOR = 8'b01010100;
localparam logic [7:0] GREEN2_COLOR = 8'b00010100;
localparam logic [7:0] TEAL_COLOR = 8'b00010000;
localparam logic [7:0] RED_COLOR = 8'b11100000;






logic [7:0][0:42][7:0] object_colors = {
{GREEN_COLOR,
 GREEN2_COLOR,
 TEAL_COLOR,
 TEAL_COLOR,
 GREEN2_COLOR,
 GREEN_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA2_COLOR,
 SEA2_COLOR,
 SEA2_COLOR},
{GREEN_COLOR,
 GREEN2_COLOR,
 GREEN2_COLOR,
 GREEN_COLOR,
 GREEN2_COLOR,
 GREEN_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA2_COLOR,
 SEA2_COLOR,
 SEA2_COLOR},
{GREEN2_COLOR,
 GREEN_COLOR,
 GREEN_COLOR,
 GREEN2_COLOR,
 GREEN_COLOR,
 GREEN2_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 WHITE_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA2_COLOR,
 SEA2_COLOR,
 SEA2_COLOR},
 {GREEN2_COLOR,
 GREEN_COLOR,
 TEAL_COLOR,
 TEAL_COLOR,
 GREEN_COLOR,
 GREEN2_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 WHITE_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA2_COLOR,
 SEA2_COLOR,
 SEA2_COLOR},
{GREEN2_COLOR,
 GREEN2_COLOR,
 GREEN_COLOR,
 GREEN_COLOR,
 GREEN2_COLOR,
 GREEN2_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 WHITE_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA2_COLOR,
 SEA2_COLOR,
 SEA2_COLOR},
 {GREEN2_COLOR,
 GREEN2_COLOR,
 GREEN_COLOR,
 GREEN_COLOR,
 GREEN2_COLOR,
 GREEN2_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 WHITE_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA2_COLOR,
 SEA2_COLOR,
 SEA2_COLOR},
{GREEN_COLOR,
 GREEN2_COLOR,
 GREEN_COLOR,
 GREEN2_COLOR,
 GREEN_COLOR,
 GREEN2_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA2_COLOR,
 SEA2_COLOR,
 SEA2_COLOR},
{GREEN_COLOR,
 GREEN2_COLOR,
 GREEN_COLOR,
 GREEN2_COLOR,
 GREEN_COLOR,
 GREEN2_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 DARK_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 LIGHT_GRAY_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SAND_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA_COLOR,
 SEA2_COLOR,
 SEA2_COLOR,
 SEA2_COLOR}
};


 
 
 
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
				BG_RGB <= BLACK_COLOR;
	end 
	else begin
	// default 
		BG_RGB <= BLACK_COLOR;
		boardersDrawReq = 0;
		 if (startOfFrame)begin
				case(speed)
					2'd1: object_colors <= {object_colors[6:0],object_colors[7]};
					2'd2: object_colors <= {object_colors[5:0],object_colors[7:6]};
					default:object_colors <= object_colors;
				endcase
			end 
		if(InsideRectangle)begin
			boardersDrawReq = 1;
			BG_RGB <= object_colors[(pixelY / 8) % 8][(pixelX/8)];
			end
		 end
end


/* logic drawingRequest;
assign drawingRequest = (BG_RGB != BLACK_COLOR ) ? 1'b1 : 1'b0 ; */
endmodule
